module judgeLess(out, i);
	input i;
	output out;
	
	and(out, i, 1'b1);

endmodule
